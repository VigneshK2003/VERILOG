module odd_parity(input a,b,c,p, output y);
	assign y = ~(a^b^c^p); 
endmodule
