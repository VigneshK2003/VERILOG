module b_to_e( input[3:0]b , output[3:0]e );
    assign e = b + 4'b0011;
endmodule

     
